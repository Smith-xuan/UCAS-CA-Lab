    `define BR_DATA_WD           34
    `define FS_TO_DS_DATA_WD     64
    `define DS_TO_ES_DATA_WD     165
    `define ES_TO_MS_DATA_WD     76
    `define MS_TO_WS_DATA_WD     70
    `define WS_TO_RF_DATA_WD     41
    `define ES_FWD_BLK_DATA_WD   42
    `define MS_FWD_BLK_DATA_WD   41