    `define BR_DATA_WD           34
    `define FS_TO_DS_DATA_WD     65
    `define DS_TO_ES_DATA_WD     192
    `define ES_TO_MS_DATA_WD     235
    `define MS_TO_WS_DATA_WD     226
    `define WS_TO_RF_DATA_WD     41
    `define ES_FWD_BLK_DATA_WD   42
    `define MS_FWD_BLK_DATA_WD   42
    `define WS_CSR_BLK_DATA_WD   15
    `define MS_CSR_BLK_DATA_WD   15 
    `define ES_CSR_BLK_DATA_WD   15 

    `define CSR_CRMD    13'h0000
    `define CSR_PRMD    13'h0001
    `define CSR_ECFG    13'h0004
    `define CSR_ESTAT   13'h0005
    `define CSR_ERA     13'h0006
    `define CSR_BADV    13'h0007
    `define CSR_EENTRY  13'h000c
    `define CSR_SAVE0   13'h0030
    `define CSR_SAVE1   13'h0031
    `define CSR_SAVE2   13'h0032
    `define CSR_SAVE3   13'h0033
    `define CSR_TID     13'h0040
    `define CSR_TCFG    13'h0041
    `define CSR_TVAL    13'h0042
    `define CSR_TICLR   13'h0044
    `define CSR_CRMD_PLV 1:0
    `define CSR_CRMD_PIE 2
    `define CSR_CRMD_DA 3
    `define CSR_PRMD_PPLV 1:0
    `define CSR_PRMD_PIE 2
    `define CSR_ECFG_LIE 12:0
    `define CSR_ESTAT_IS10 1:0
    `define CSR_ERA_PC 31:0
    `define ECODE_ADE 6'b001000
    `define ECODE_ALE 6'b001001
    `define ESUBCODE_ADEF 9'b0
    `define CSR_EENTRY_VA 31:6
    `define CSR_SAVE_DATA 31:0
    `define CSR_TID_TID 31:0
    `define CSR_TCFG_EN 0
    `define CSR_TCFG_PERIOD 1
    `define CSR_TCFG_INITV 31:2
    `define CSR_TICLR_CLR 0
